package bt_top;

parameter int ADDR_WIDTH = 8;
parameter int BURST_LEN = 15;
parameter int DATA_WIDTH = 8;

endpackage



package sram_pkg;

parameter int ADDR_WIDTH = 8;
parameter int DATA_WIDTH = 8;

endpackage //sram_pkg